LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY UART_DATA IS
	PORT(
		CLOCK    : IN    STD_LOGIC;
		RESETN   : IN    STD_LOGIC;
		CS		 : IN	 STD_LOGIC;
		UART_STB : IN    STD_LOGIC;
		IO_DATA  : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END UART_DATA;


ARCHITECTURE a OF UART_DATA IS
	SIGNAL IO_OUT : STD_LOGIC;
	SIGNAL OUTDATA : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
	-- Use LPM function to drive I/O bus
	IO_BUS: LPM_BUSTRI
	GENERIC MAP (
		lpm_width => 16
	)
	PORT MAP (
		data     => OUTDATA,
		enabledt => IO_OUT,
		tridata  => IO_DATA
	);
	
	IO_OUT <= CS;

	PROCESS (CLOCK, RESETN)

	BEGIN
		IF (RESETN = '0') THEN          -- Active low, asynchronous reset
			OUTDATA <= x"0000";
		ELSIF (RISING_EDGE(CLOCK)) THEN
			OUTDATA <= (x"000" & "000" & UART_STB);
		END IF;
	END PROCESS;
END a;